Sin fondo